module key2asc(
    input [7:0] keybuffer,
    output reg [11:0] asci 

);
    MuxKeyWithDefault#(67, 8, 12) key2ascMux(.out(asci), .key(keybuffer), .default_out(12'b1111_1111_1111), .lut({
	8'h1C, 12'h065,
	8'h32, 12'h066,
    8'h21, 12'h067,
    8'h23, 12'h068,
    8'h24, 12'h069,
    8'h2B, 12'h070,
    8'h34, 12'h071,
    8'h33, 12'h072,
    8'h43, 12'h073,
    8'h3B, 12'h074,
    8'h42, 12'h075,
    8'h4B, 12'h076,
    8'h3A, 12'h077,
    8'h31, 12'h078,
    8'h44, 12'h079,
    8'h4D, 12'h080,
    8'h15, 12'h081,
    8'h2D, 12'h082,
    8'h1B, 12'h083,
    8'h2C, 12'h084,
    8'h3C, 12'h085,
    8'h2A, 12'h086,
    8'h1D, 12'h087,
    8'h22, 12'h088,
    8'h35, 12'h089,
    8'h1A, 12'h090,
    8'h45, 12'h048,
    8'h16, 12'h049,
    8'h1E, 12'h050,
    8'h26, 12'h051,
    8'h25, 12'h052,
    8'h2E, 12'h053,
    8'h36, 12'h054,
    8'h3D, 12'h055,
    8'h3E, 12'h056,
    8'h05, 12'h112,
    8'h06, 12'h113,
    8'h04, 12'h114,
    8'h0C, 12'h115,
    8'h03, 12'h116,
    8'h0B, 12'h117,
    8'h83, 12'h118,
    8'h0A, 12'h119,
    8'h01, 12'h120,
    8'h09, 12'h121,
    8'h78, 12'h122,
    8'h07, 12'h123,
    8'h66, 12'h008,
    8'h0D, 12'h009,
    8'h5A, 12'h013,
    8'h12, 12'h016,
    8'h14, 12'h017,
    8'h11, 12'h018,
    8'h58, 12'h020,
    8'h76, 12'h027,
    8'h29, 12'h032,
    8'h4C, 12'h186,
    8'h55, 12'h187,
    8'h41, 12'h188,
    8'h4E, 12'h189,
    8'h49, 12'h190,
    8'h4A, 12'h191,
    8'h0E, 12'h192,
    8'h54, 12'h219,
    8'h5B, 12'h221,
    8'h5D, 12'h220,
    8'h52, 12'h222
	}));
endmodule