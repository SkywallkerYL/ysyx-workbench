module ysyx_22050550_EXU (
    
);
    
endmodule